package cpu_package is

constant DATA_WIDTH_C			: positive := 32;
constant NUM_REGS_C				: positive := 32;
constant NUM_ALU_CTRL_C			: positive := 4;

end package;